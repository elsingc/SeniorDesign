`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:07:06 12/15/2013 
// Design Name: 
// Module Name:    Accelerometer_Controller 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Accelerometer_Controller(
	output [19:0] x_accl,
	output [19:0] y_accl,
	output [19:0] z_accl,
	output ena,
	output [7:0] data_wr,
	output [7:0] data_rd,
	input busy,
	output new,
	input rst,
	input clk
    );


endmodule
