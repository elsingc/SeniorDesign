`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:15:09 12/15/2013 
// Design Name: 
// Module Name:    Camera_Digitizer 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Camera_Digitizer(
	input busy,
	input block,
	input new_data,
	input [7:0] data,
	input dtr,
	input vsync,
	input href,
	input pclk,
	input [7:0] ybus,
	input rst,
	input clk
    );


endmodule
