`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:10:09 12/15/2013 
// Design Name: 
// Module Name:    Analog_Controller 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Analog_Controller(
	output [7:0] ch0,
	output [7:0] ch1,
	output [7:0] ch4,
	output [7:0] ch5,
	output [7:0] ch6,
	output [7:0] ch7,
	output [7:0] ch8,
	output [7:0] ch9,
	output [7:0] channel,
	input new_sample,
	input [7:0] sample,
	input [7:0] sample_channel,
	input rst,
	input clk
    );


endmodule
